module decoder38_15 (i_sel, i_opt, o_y);
    input [2:0] i_sel;
    input i_opt;
    output [7:0] o_y;
    reg [7:0] r_y;
    
endmodule
